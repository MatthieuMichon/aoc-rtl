`timescale 1ns/1ps
`default_nettype none

module user_logic (
    input wire tck,
    input wire tdi,
    output logic tdo,
    input wire test_logic_reset,
    input wire run_test_idle,
    input wire ir_is_user,
    input wire capture_dr,
    input wire shift_dr,
    input wire update_dr
);

localparam int BYTE_WIDTH = $bits(byte);
// From design space exploration
localparam int RESULT_WIDTH = 16;
parameter int DEVICE_CHARS = 3;
parameter int DEVICE_BIN_BITS = 5;
parameter int DEVICE_WIDTH = DEVICE_CHARS*DEVICE_BIN_BITS;
parameter int MAX_NODES = 1024;
parameter int NODE_WIDTH = $clog2(MAX_NODES);

typedef logic [NODE_WIDTH-1:0] node_t;

logic inbound_valid;
logic [BYTE_WIDTH-1:0] inbound_data;

tap_decoder #(.DATA_WIDTH(BYTE_WIDTH)) tap_decoder_i (
    // TAP signals
        .tck(tck),
        .tdi(tdi),
        .test_logic_reset(test_logic_reset),
        .ir_is_user(ir_is_user),
        .shift_dr(shift_dr),
        .update_dr(update_dr),
    // Decoded signals
        .valid(inbound_valid),
        .data(inbound_data)
);

logic decoding_done_str;
logic edge_str_valid;
logic src_node_str_valid;
logic [DEVICE_WIDTH-1:0] src_node_str;
logic [DEVICE_WIDTH-1:0] dst_node_str;

input_decoder input_decoder_i (
    .clk(tck),
    // Inbound Byte Stream
        .byte_valid(inbound_valid),
        .byte_data(inbound_data),
    // Decoded signals
        .decoding_done(decoding_done_str),
        .edge_valid(edge_str_valid),
        .src_node_valid(src_node_str_valid),
        .src_node(src_node_str),
        .dst_node(dst_node_str)
);

logic decoding_done_idx;
logic edge_idx_valid;
logic src_node_idx_valid;
node_t src_node_idx;
node_t dst_node_idx;
node_t node_idx_cnt;
node_t start_node_idx;
node_t end_node_idx;
logic start_end_nodes_valid;

node_id_mapper node_id_mapper_i (
    .clk(tck),
    // Node with Random Identifier
        .decoding_done_str(decoding_done_str),
        .edge_str_valid(edge_str_valid),
        .src_node_str_valid(src_node_str_valid),
        .src_node_str(src_node_str),
        .dst_node_str(dst_node_str),
    // Node with Indexed Identifier
        .decoding_done_idx(decoding_done_idx),
        .edge_idx_valid(edge_idx_valid),
        .src_node_idx_valid(src_node_idx_valid),
        .src_node_idx(src_node_idx),
        .dst_node_idx(dst_node_idx),
        .node_idx_cnt(node_idx_cnt),
    // Static Start and End Nodes
        .start_node_idx(start_node_idx),
        .end_node_idx(end_node_idx),
        .start_end_nodes_valid(start_end_nodes_valid)
);

logic query_ready;
logic query_valid;
node_t query_data;
logic reply_ready;
logic reply_valid;
logic reply_last;
node_t reply_data;
logic reply_no_edges_found;

adjacency_map adjacency_map_i(
    .clk(tck),
    // Connection Entries
        .decoding_done(decoding_done_idx),
        .edge_valid(edge_idx_valid),
        .src_node_valid(src_node_idx_valid),
        .src_node(src_node_idx),
        .dst_node(dst_node_idx),
    // Query/Reply Interface
        .query_ready(query_ready),
        .query_valid(query_valid),
        .query_data(query_data),
        .reply_ready(reply_ready),
        .reply_valid(reply_valid),
        .reply_last(reply_last),
        .reply_data(reply_data),
        .reply_no_edges_found(reply_no_edges_found)
);

node_t indeg_node;
logic indeg_dec;
node_t indeg_degree;

indegree_list indegree_list_i (
    .clk(tck),
    // Connection Entries
        .edge_valid(edge_idx_valid),
        .dst_node(dst_node_idx),
    // Update Interface
        .node_sel(indeg_node),
        .decrement_degree(indeg_dec),
        .node_degree(indeg_degree) // degree after decrement
);

logic sorted_done;
logic sorted_valid;
node_t sorted_node;

topological_sort topological_sort_i (
    .clk(tck),
    // Connection Entries
        .decoding_done(decoding_done_idx),
        .node_idx_cnt(node_idx_cnt),
    // Indegree List Interface
        .indeg_node(indeg_node),
        .indeg_dec(indeg_dec),
        .indeg_degree(indeg_degree), // degree after decrement
    // Query/Reply Interface
        .query_ready(query_ready),
        .query_valid(query_valid),
        .query_data(query_data),
        .reply_ready(reply_ready),
        .reply_valid(reply_valid),
        .reply_last(reply_last),
        .reply_data(reply_data),
        .reply_no_edges_found(reply_no_edges_found),
    // Sorted Nodes
        .sorted_done(sorted_done),
        .sorted_valid(sorted_valid),
        .sorted_node(sorted_node)
);

logic trimed_done;
logic trimed_valid;
node_t trimed_node;

node_list_trim node_list_trim_i (
    .clk(tck),
    // Node with Indexed Identifier
        .start_node_idx(start_node_idx),
        .end_node_idx(end_node_idx),
        .start_end_nodes_valid(start_end_nodes_valid),
    // Sorted Nodes
        .sorted_done(sorted_done),
        .sorted_valid(sorted_valid),
        .sorted_node(sorted_node),
    // Trimed Sorted Nodes
        .trimed_done(trimed_done),
        .trimed_valid(trimed_valid),
        .trimed_node(trimed_node)
);

// logic debug_valid____;
// logic [16-1:0] debug_cnt____;

// always_ff @(posedge tck) begin
//     if (trimed_valid) begin
//         debug_cnt____ <= debug_cnt____ + 1;
//     end
// end
// assign debug_valid____ = trimed_done;

logic outbound_valid;
logic [RESULT_WIDTH-1:0] outbound_data;

node_path_counter node_path_counter_i (
    .clk(tck),
    // Adjacency Nodes Entries
        .decoding_done(decoding_done_idx),
        .edge_valid(edge_idx_valid),
        .src_node_valid(src_node_idx_valid),
        .src_node(src_node_idx),
        .dst_node(dst_node_idx),
    // Matching Indexes for Start/End Nodes
        .start_node_idx(start_node_idx),
        .end_node_idx(end_node_idx),
        .start_end_nodes_valid(start_end_nodes_valid),
    // Sorted Nodes
        .trimed_done(trimed_done),
        .trimed_valid(trimed_valid),
        .trimed_node(trimed_node),
    // Path Count
        .path_count_valid(outbound_valid),
        .path_count_value(outbound_data)
);

tap_encoder #(.DATA_WIDTH(RESULT_WIDTH)) tap_encoder_i (
    // TAP signals
        .tck(tck),
        .tdo(tdo),
        .test_logic_reset(test_logic_reset),
        .ir_is_user(ir_is_user),
        .capture_dr(capture_dr),
        .shift_dr(shift_dr),
    // Encoded signals
        .valid(outbound_valid),
        .data(outbound_data)
);

wire _unused_ok = 1'b0 && &{1'b0,
    start_node_idx,
    trimed_done,
    trimed_node,
    sorted_node,
    src_node_idx_valid,
    src_node_idx,
    dst_node_idx,
    node_idx_cnt,
    start_node_idx,
    end_node_idx,
    start_end_nodes_valid,
    src_node_str_valid,
    src_node_str,
    dst_node_str,
    edge_str_valid,
    run_test_idle,  // To be fixed
    1'b0};

endmodule
`default_nettype wire
